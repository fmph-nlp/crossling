<s snum=1> Detta åtagande är viktigt , med tanke på att kommissionen är det organ som enligt fördragen har ensam initiativrätt , och det utgör därför grunden till parlamentets politiska och lagstiftande verksamhet de kommande fem åren . </s>
<s snum=2> ( Applåder ) Det är sista gången vi tar hänsyn till att ni glömt korten . </s>
<s snum=3> Jag kommer ju , precis_som min kollega Rack , från ett transitland , där denna fråga spelar en särskild roll . </s>
<s snum=4> Vid en av de större olyckor som inträffat på senare tid , var inte det transporterade godset farligt i sig . </s>
<s snum=5> Vi vänder oss till kommissionen för att ta itu med frågor som har att göra med kompletterande medel . </s>
<s snum=6> Det är ungdomarna som försvinner , som utbildar sig och får arbete i städerna , något som påverkar landsbygden på ett negativt sätt . </s>
<s snum=7> Herr talman , herr kommissionär , värderade kolleger ! Även jag skulle vilja gratulera föredraganden och tacka henne för hennes stora och seriösa arbetsinsats . </s>
<s snum=8> Den första är den väsentliga och centrala betydelse som vi fortfarande fäster vid den ekonomiska och sociala sammanhållningen . </s>
<s snum=9> Det är själva texten jag citerat , inom citationstecken . </s>
<s snum=10> Detta kan till stor del förklaras av strukturfonderna , även_om skillnaderna mellan de fattigaste och de rikaste områdena fortfarande är avsevärda . </s>
<s snum=11> Herr talman , mina damer och herrar , kära kolleger ! Kommissionens vitbok om modernisering av de europeiska konkurrensreglerna har utlöst en intensiv och livlig debatt bland den intresserade allmänheten . </s>
<s snum=12> Reaktionerna från experter och berörda parter sträcker sig från totalt avvisande till förbehållslöst stöd . </s>
<s snum=13> Samtidigt är skillnaderna mellan staterna avsevärda och kan bedömas på olika sätt , bl.a. i procent av mervärdet och per löntagare . </s>
<s snum=14> Kommissionen måste bedriva klappjakt på illegala stöd och de stöd som verkligen blockerar den inre marknaden . </s>
<s snum=15> Jag anser att det även är den förda konkurrenspolitiken som bär ansvaret för allt detta , och jag tar fullständigt avstånd från den . </s>
<s snum=16> Men vi måste vara vaksamma när det gäller de aktörer som verkar över hela världen , som det nationella agerandet inte längre kan sätta några gränser för . </s>
<s snum=17> Fyrtio år senare dyker detta förslag nu upp igen , och det kommer - det är jag säker på - att ge utrymme för kartellbildningar till nackdel för konsumenterna i Europa . </s>
<s snum=18> Jag måste dock säga att min grupp tyvärr inte kommer att rösta enhälligt för ert betänkande . </s>
<s snum=19> Med den_här texten rör vi oss verkligen i utkanten av vad_som är möjligt , eftersom vi anser att det finns frågor som måste lösas och att det är viktigt att bedrägerierna inom gemenskapen stoppas , att de stryps . </s>
<s snum=20> I egenskap av ledamot av Europaparlamentet för Leinsters valkrets har jag alltid hävdat behovet av att förverkliga lokala initiativ som stöds av nationella EU-fonder . </s>
<s snum=21> Under dessa tragiska omständigheter tror jag att det vore en missuppfattning och en skam om vi talade med flera olika röster , principiellt sett . </s>
<s snum=22> Jag vill be staterna att gripa tag i det tillfället : detta program måste fungera fullt ut . </s>
<s snum=23> Denna situation skapas inte genom myndighetens blotta tillkomst utan kommer att framträda efter hand i takt med att självförtroendet stiger inom myndigheten själv . </s>
<s snum=24> Upprättandet av den positiva listan är en av de frågor som behandlas i bilagan som har ett datum åsatt , år 2002 faktiskt . </s>
<s snum=25> Europeiska kommissionen har övervakat konfliktens miljökonsekvenser från det att Natoaktionen inleddes . </s>
<s snum=26> Jag kan inte svara på den frågan . </s>
<s snum=27> Frågan är nu vad kommissionen kan göra för att på ett mer konkret sätt stödja Hans Helighet Dalai Lama och hans förslag till en fredlig lösning av Tibet-frågan ? </s>
<s snum=28> Detta begränsade utbildningsmoment har dock strukits från alla introduktionskurser som har ägt rum under senare tid . </s>
<s snum=29> Avsatta medel för de icke-statliga organisationernas program i Tadzjikistan uppgick till 7,42 miljoner euro 1998 och 1999 . </s>
<s snum=30> Jag är mycket mån om att vi stärker våra relationer med dem . </s>
<s snum=31> Vid Europeiska rådets möte i Lissabon görs ett nytt försök att ta itu med frågan om den sociala utslagningen , den sociala utslagningens samband med informationssamhället , med den ekonomiska politiken och med reformerna . </s>
<s snum=32> Det är ett utmärkt betänkande och vi bör alla gratulera henne till det . </s>
<s snum=33> Även här vill jag försäkra att ni där berör en av de reformer som kommissionen syftar till . </s>
<s snum=34> Detta är väsentligt för ett verkställande organ som skall vara redovisningsskyldigt , inte_bara inför detta parlament , utan mer generellt inför den europeiska allmänheten . </s>
<s snum=35> En varaktig fred i det_här området kan förverkligas först genom ett avtal i vilket säkerheten för de israeliska gränserna och Syriens integritet kan garanteras . </s>
<s snum=36> Herr talman , kommissionär Patten , kära kolleger ! </s>
<s snum=37> Men jag vill påminna ordförande Prodi om att han i utnämningsdebatten talade om kommissionen som en europeisk regering . </s>
<s snum=38> Men vi var också upprörda över vänsterns överseende med tyranniet , terrorn och övergreppen i f.d. Sovjetunionen . </s>
<s snum=39> I första hand värdena och principerna om frihet , demokrati och respekt för de mänskliga rättigheterna . </s>
<s snum=40> Har ni någon gång frågat er om vi inte också är ansvariga för den fortsatta utvecklingen av det politiska läget i Österrike , om vi här sätter oss till doms över detta ? </s>
<s snum=41> Men det är sant att det krävs inte uppbackning av en stor majoritet av det vetenskapliga samfundet för att kunna använda försiktighetsprincipen . </s>
<s snum=42> Tack , fru kommissionär . </s>
<s snum=43> Vi skall inte längre oroa oss över att dagordningen för regeringskonferensen skall bli begränsad . </s>
<s snum=44> Det vi behöver är synliga rättigheter för var_och_en , stadgan om de grundläggande rättigheterna måste blir bindande rätt för alla människor som bor i unionen , för alla dess medborgare . </s>
<s snum=45> Fördragets artikel 56 , som förbjuder varje ingrepp i den fria rörligheten för kapitalet , valutaspekulationen , måste tas bort så att den skadliga valutaspekulationen kan hejdas genom politisk kontroll . </s>
<s snum=46> Det kan dessutom fastslås att av 19 departement har redan 4 en administrativ ledning , vilket också är ett framsteg jämfört med vad vi tidigare haft där . </s>
<s snum=47> Detta är händelser och situationer som vi inte kan acceptera . </s>
<s snum=48> Jo , i enkla ekonomiska termer främjar europeisk kultur verkligt välstånd . </s>
<s snum=49> Jag anser det inte nödvändigt att veteranbilar skall utgöra en_del av direktivet . </s>
<s snum=50> Det är mitt huvudsakliga bekymmer på det området . </s>
<s snum=51> I så måtto föreslår jag att en fond för de gamla fordonen bildas , ur vilken återvinningskostnaderna för de uttjänta fordonen sedan betalas så att principen om kostnadsbefrielse säkras . </s>
<s snum=52> Vi diskuterar denna fråga i ett annat forum i parlamentet . </s>
<s snum=53> Det finansieras via en fond som nybilsköparna betalar in till . </s>
<s snum=54> Jag anser att detta är en graverande brist som i princip inte heller passar vårt rättssystem . </s>
<s snum=55> Valet till Europaparlamentet 1999 visade med all tydlighet att medborgarna inte följer med i tankegångarna om ett allt mer Brysselfederalistiskt EU . </s>
<s snum=56> Jag har noterat era budskap i frågan och jag tror att Banotti har ett svar till er . </s>
<s snum=57> Jag anser att frågan är så viktig att vi bör följa den , men inte att vi skall lösa den med hjälp av förfarandet för brådskande ärenden . </s>
<s snum=58> Det är denna typ av bra åtgärder som vi också vill skall utvidgas till hela EU när det rör kommunikation och offentlighet . </s>
<s snum=59> Nu tycks också de stödåtgärder som anförs i bilaga II till programinriktning A vara lovande i detta hänseende . </s>
<s snum=60> Vissa områden i Europeiska unionen är ekonomiskt sett mycket starka och överskrider mycket tydligt den genomsnittliga inkomsten per_capita . </s>
<s snum=61> De gröna kan därför inte räkna med vårt stöd för ändringsförslag 2 , vilket de inte heller fick under utskottssammanträdet . </s>
<s snum=62> Att vara solidarisk med Östeuropa är nog bra , men det räcker inte . </s>
<s snum=63> Vi beklagar , precis_som föredraganden , att kapitel IIIA har tagits bort . </s>
<s snum=64> Till_sist några ord om Interreg . </s>
<s snum=65> Det var mitt första svar på frågan om tröskeln . </s>
<s snum=66> Dessa är våra stora handlingslinjer för de kommande fem åren . </s>
<s snum=67> Det är dags att fundera på , och sedan förverkliga , en europeisk räddningstjänst . </s>
<s snum=68> Men vi säger också att vi vill försvara detta europeiska samhälle av tolerans , och därför är en gemensam utrikes - , säkerhets - och försvarspolitik så viktig . </s>
<s snum=69> Vi får inte låta kritikerna av europeisk integration hävda , som de för_närvarande gör med visst berättigande enligt vad vi just har hört av Bonde , att ökningen av EU : s ansvarsområden endast går åt ett håll . </s>
<s snum=70> Europa som är så demokratiskt , som är så progressivt , tiger och tar inte på sig dessa tragiska problem , under tiden som halva Afrika dör i aids och andra sjukdomar . </s>
<s snum=71> En union enbart som ett geostrategiskt koncept har inte någon framtid , lika litet som en union som enbart är en frihandelszon . </s>
<s snum=72> Herr talman ! Enligt Europeiska liberala och demokratiska partiets grupp är kommissionens och hela unionens viktigaste uppgift under de närmaste åren att genomföra utvidgningen med framgång . </s>
<s snum=73> Det nya Europa får inte_bara utvecklas på bredden utan_även på djupet , genom att omsätta våra värden i praktiken och genom ett demokratiskt byggande av en äkta gemenskap . </s>
<s snum=74> De regeringar som stöder er av slapphet eller av ideologiska skäl är det också . </s>
<s snum=75> Vi är och kommer att förbli bland dem som bekämpar en europeistisk diktatur och vi uppmanar alla Europas folk att gå med i motståndet mot era ohyggliga förslag . </s>
<s snum=76> Vilken bild får då en intresserad allmänhet och resten av världen av detta femårsprogram ? </s>
<s snum=77> Med instämmande i vad mina partivänner har sagt och med gillande av grundtonen i ert dokument vill jag rikta uppmärksamheten på två brister , som måste korrigeras i det kommande arbetet . </s>
<s snum=78> Alla vet att livskvalitet , full sysselsättning och bättre sysselsättning är beroende av en hållbar ekonomisk tillväxt . </s>
<s snum=79> Nästan 40 procent av företagen i denna undersökning meddelar att de fortfarande har extra omkostnader för att göra produkter eller tjänster förenliga med nationella specifikationer . </s>
<s snum=80> Det skulle vara tragiskt om deras ansträngningar skulle undergrävas på_grund_av brister i EU : s lagstiftning . </s>
<s snum=81> Vi skall granska i vilken omfattning vi kan skapa en liksidig triangelformad politik där man kombinerar ekonomisk politik , sysselsättningspolitik och socialpolitik . </s>
<s snum=82> Herr talman ! Även jag vill ta upp en ordningsfråga . </s>
<s snum=83> Personligen anser jag att det är inget mindre än skandal att vi har ledamöter i detta parlament som angriper demonstrationen hellre än att söka lösningen på problemet , vilket är rimliga arbetsförhållanden , rimlig lön och rimliga arbetstider . </s>
<s snum=84> Vi kan aldrig tillräckligt påminna om de svårigheter som fanns förr i tiden i de områden vid gränserna , på land eller till havs , som hade delats ekonomiskt , socialt och kulturellt . </s>
<s snum=85> Detta framgår av det faktum att jordbruksinkomsterna och sysselsättningen har minskat mycket hastigt i de områden där dessa initiativ har tillämpats , vilket lett till allt snabbare avfolkning av dessa områden . Grekland är ett betecknande exempel . </s>
<s snum=86> Kommissionen föreslog att införa en rättslig grund från och med oktober 1999 i direktiv 70 / 524 / EEG för att ersätta tillstånden . </s>
<s snum=87> Det får ändå inte vara så att ni undantar kosmetika , farmaceutika och andra produkter med motiveringen att det inte kan uppstå några skador eller att det inte är farligt . </s>
<s snum=88> I det aktuella förslaget har jag föreslagit att man skall stryka alla nu gällande gemenskapsbestämmelser om skrapie hos får och getter och att införliva dem i ramförslaget om en förordning . </s>
<s snum=89> Många direktiv har antagits och kommissionens vilja är för_övrigt att lyckas med att göra dem läsbarare , mer överensstämmande sinsemellan samt förse dem med tydligare mål . </s>
<s snum=90> Vi måste försöka få till stånd ett medlingsförfarande . </s>
<s snum=91> För ungefär sju år sedan verkade det också som_om den europeiska vattenpolitiken skulle offras på subsidiaritetsaltaret . </s>
<s snum=92> Vi har inte råd att vänta . </s>
<s snum=93> Herr talman ! Jag uppskattar Barniers löfte att gå ut till regionerna , både för att förklara och för att lyssna till vad medborgarna har att säga . </s>
<s snum=94> Utvecklingen går långsamt på_grund_av de spända förbindelserna mellan de etniska grupperna i denna delade stad . </s>
<s snum=95> Jag var i Mitrovica för några månader sedan och såg själv situationen där . </s>
<s snum=96> Föregående fråga föranledde oss att tala om valen . </s>
<s snum=97> Får jag be att få tacka herr Andersson för fortsättningen på hans första fråga och den frågan vill jag svara på så_här . </s>
<s snum=98> Om jag förstått det rätt så har Posselt börjat peka på skatteaspekterna av den_här frågan . </s>
<s snum=99> Även_om vi kommer fram_till vem_som beslutar om sådana ingrepp , anser jag att vi behöver gemensamma och mycket stränga regler . </s>
<s snum=100> Detta reflekteras också i flera av parlamentets ändringsförslag . </s>
<s snum=101> Nitratdirektivet kommer därför inte att påverkas av detta ramdirektiv . </s>
<s snum=102> I ändringsförslag 71 tas inte hänsyn till årtidsvariationer och årliga förändringar i grundvattennivån . </s>
<s snum=103> Herr talman ! Först av allt vill jag gratulera Lienemann till den starka känsla för miljöfrågorna som märks i de två betänkanden vi diskuterar i kväll . </s>
<s snum=104> Verkligheten är helt annorlunda . </s>
<s snum=105> Och detta är det paradoxala . </s>
<s snum=106> Här omfattas även personer från tredje land och statslösa personer . </s>
<s snum=107> Den allmännyttiga politiska samstämmigheten är därför ett ansvar för kommissionen som helhet , för rådet och för Europaparlamentet . </s>
<s snum=108> Jag vill särskilt framhålla att det verkar som_om vi börjar få ett nytt sätt att se på de_här frågorna , främst när det gäller handel , något som var välbehövligt . </s>
<s snum=109> På samma sätt som för styrkeförhållandena som studeras inom den elementära fysiken är det ingen mening med att införa politikområden som motverkar varandra . </s>
<s snum=110> Den skulle även behöva snabbare kontrakts - och tillämpningsförfaranden samt en utökad flerårig budgetpost och en kraftigt förbättrad förvaltning av sina program . </s>
<s snum=111> Alla känner vi till rapporterna från Amnesty International . </s>
<s snum=112> OMRÖSTNING ( fortsättning ) </s>
<s snum=113> Debatterna om försiktighetsprincipen , spårbarhet , ansvar och öppenhet har förmått Europeiska kommissionen att presentera en vitbok om livsmedelssäkerhet . </s>
<s snum=114> Enligt min åsikt är det felaktigt att använda ett så trubbigt verktyg som en gemensam europeisk avgift i denna fråga . </s>
<s snum=115> Vi har blivit vittnen till hur ett betänkande som värnar om Europas vattenkvalitet förvandlas till ett instrument i ett handelskrig . </s>
<s snum=116> FN : s nästa session om mänskliga rättigheter ( fortsättning ) </s>
<s snum=117> Hur genomför vi det som föreskrivs i fördragen i alla dessa ord om utvecklingsbiståndsprogram ? </s>
<s snum=118> Finns det möjlighet att avstänga honom från sin befattning till det att den rättsliga undersökningen slutförts ? </s>
<s snum=119> Ni antydde det nyss , här står vi inför en katastrof , och ingenting görs . </s>
<s snum=120> Kosovoproblemet är känt ; där finns världssamfundet närvarande i stor omfattning . </s>
<s snum=121> Det har även tagits ett litet steg , som hör samman med det partiella upphävandet nyligen av embargot mot Jugoslavien , vilket beslutades av våra 15 regeringar . </s>
<s snum=122> Det är viktigt att i tid ha ett straffrättsligt skydd i alla länder som ser någorlunda likadant ut . </s>
<s snum=123> Tack även till dem som har bidragit till en snabb hantering i frågan ; jag tänker särskilt på PSE-gruppen . </s>
<s snum=124> Varje stat måste därmed se till att effektiva straffpåföljder införs , påföljder som skall vara lämpliga och avskräckande för de brott som förutses i förslaget till rambeslut . </s>
<s snum=125> Vi har kommit fram_till att så inte är fallet , men med tanke på hur viktigt ämnet är har vi ändå enats om att acceptera förfarandet . </s>
<s snum=126> Protokollet från i_går har delats ut . </s>
<s snum=127> Några av ändringsförslagen går dock för långt i att begränsa användandet av OTC-derivat . </s>
<s snum=128> Master - / Feeder-fonder står följaktligen i motsatsställning till avsikten i direktivet och har av den anledningen helt korrekt avvisats av utskottet för ekonomi och valutafrågor . </s>
<s snum=129> Även_om vi i utskottet för ekonomi och valutafrågor i mycket var eniga om målsättningarna i lagstiftningsreformen var inte utskottsbehandlingen bland de allra lättaste . </s>
<s snum=130> Detta kumulativa villkor är väsentligt , eftersom straffrättens legalitetsprincip " nulla poena sine lege " enligt min uppfattning bör respekteras . </s>
<s snum=131> Förutom det så har Europeiska rådet i Tammerfors redan visat i vilken riktning vi , i kommissionen , borde gå . </s>
<s snum=132> Men nu vill Prodi-kommissionen göra om EU för att aspirera på posten som internationell ledare vid sidan av Förenta_staterna , samtidigt_som vi skall tävla och konkurrera med dem . </s>
<s snum=133> Vi är väl medvetna om den aktuella ekonomiska bakgrunden , eftersom omstruktureringarna syftar till att rationalisera förvaltningen av företagen . </s>
<s snum=134> Vad beträffar kan vi för_närvarande se ett antal stora fusioner som kommer till stånd mellan företag som kommer från den anglosaxiska traditionen och företag som snarare kommer från Rhenlandets tradition . </s>
<s snum=135> Alltid när ett allvarligt socialt problem uppträder finns det en politisk bakgrund : detta är vår åsikt angående de olyckliga händelserna nyligen i El Ejido . </s>
<s snum=136> Det som hände i El Ejido avslöjar otillåtliga rasistiska och främlingsfientliga metoder i dagens Europa . </s>
<s snum=137> Deras enda brott består av att de kritiserat det som människorättsorganisationer sedan_länge har klagat på , nämligen den storskaliga korruptionen och de hundratals miljoner dollar , utbetalade av oljebolagen till den angolanska regeringen , som försvunnit . </s>
<s snum=138> Ursprungsbefolkningen i USA - Dineh </s>
<s snum=139> De är bara några få , men deras motståndare är en mycket mäktig ekonomisk faktor . </s>
<s snum=140> Det blev jag övertygad om i Sarajevo när jag fick agera för att förhandla med konfliktens parter om regelbundna utväxlingar av fångar , som följde på varje eld-upphör-avtal , tyvärr aldrig särskilt varaktiga . </s>
<s snum=141> Frågan är alltså : vilka krav måste vi eventuellt ställa på ett monopol eller en_del av en tjänst som domineras av ett monopol ? </s>
<s snum=142> Avregleringen har alltså avlägsnat många parasiter inom många områden och gjort det möjligt för många att få en högre levnadsstandard . </s>
<s snum=143> Det talades om landsbygden , om glesbefolkade områden . </s>
<s snum=144> I en värld av nätverk är posten det mest demokratiska nätverket . </s>
<s snum=145> Vi har en mycket högt kvalificerad personal med en kompetens som det är svårt - kanske omöjligt - att hitta i de enskilda ländernas byråkratier , just på_grund_av hur personalen rekryteras och de urvalskriterier som tillämpas . </s>
<s snum=146> ( Kommissionären visade att han ville ha ordet senare . ) Då så , tack . </s>
<s snum=147> Man riskerar livet i Kosovo , men det är priset för friheten just nu . </s>
<s snum=148> Sedan sex månader för de ryska ledarna ett smutsigt krig av kolonialtyp , på_grund_av simpla maktambitioner , vilket leder till en daglig dos av barbari . </s>
<s snum=149> Denna önskan infriades dock inte av Europeiska rådet vid toppmötet i Helsingfors i slutet av förra året . </s>
<s snum=150> Min andra fråga är annorlunda , även_om den också har koppling till den föregående . </s>
<s snum=151> Solana kan spela en viktig roll . </s>
<s snum=152> Premiärministrar , ledamöter , bankirer , ministrar , på yrkeslivets arena , läkare , domare , piloter , militärer . </s>
<s snum=153> Problemet är att finna ändamålsenliga lösningar som medger ett större antal kvinnor på ansvarsfulla poster och därmed i beslutsfattandet . </s>
<s snum=154> Vad det rör sig om kan väl knappast uttryckas klarare än så . </s>
<s snum=155> Nu fokuserar vi i dag på hur fler kvinnor skall kunna delta i beslutsprocessen . </s>
<s snum=156> Och vi måste säga det mycket tydligt , detta sker genom ytterligare besparingar i tjänster , ytterligare tredelade system , ytterligare minskad genomsnittlig arbetstid , oavsett vilken metod vi väljer för att uppnå detta . </s>
<s snum=157> För det tredje är vi fullständigt överens om att arbetsrelationerna i Europa måste reformeras , men det betyder i klartext för oss att vi måste bevara och berika humankapitalet . </s>
<s snum=158> Vissa uppgifter är inte lämpliga , precis_som man påpekade , till_exempel sådana som handlar om beskattningen av företag . </s>
<s snum=159> Av detta landades 80 procent med snörpvad . </s>
<s snum=160> Här kan och får vi inte stå handlingsförlamade och titta på . </s>
<s snum=161> Principen att förorenaren betalar tycks oss , förutom att den är nödvändig , lämplig . </s>
<s snum=162> Den franska regeringen har lagt fram idéer och förslag för att stärka säkerheten till havs , bland_annat genom att motarbeta bekvämlighetsflagg och genomföra mycket mer omfattande kontroller . </s>
<s snum=163> Jag vill inte heller att vår muntliga fråga tas emot som ett angrepp . </s>
<s snum=164> Vi har valt att lägga ned våra röster i omröstningen om ändringsförslag 4 i Katiforisbetänkandet om Ekonomin i unionen ( 1999 ) . </s>
<s snum=165> Kan vi verkligen uppnå full sysselsättning utan att släppa lös den företagstalangen ? </s>
<s snum=166> Och Europa behöver nå upp_till en full sysselsättning . </s>
<s snum=167> Tack så mycket , herr kommissionär ! </s>
<s snum=168> Ändå fanns det i första behandlingen en_hel_del ändringsförslag och de står parlamentet helt bakom . </s>
<s snum=169> Det enda som skiljer oss åt är hur man bäst skall uppnå det . </s>
<s snum=170> Vi måste också ha klart för oss , herr kommissionsordförande , att man redan nu måste börja med dessa kriterier och detta arbete . </s>
<s snum=171> Förra månaden talade Prodi om en genomgripande decentralisering av unionens verksamhet . </s>
<s snum=172> Vi skulle inte längre sitta i utskottsrummen och titta på studenterna som bakvägen från de permanenta representationerna har de handlingar som vi inte kunde få . </s>
<s snum=173> Bättre levnadsvillkor , sysselsättning och sysselsättningens kvalitet förblir nära förbundna med vår förmåga att göra den europeiska forskningen dynamisk . </s>
<s snum=174> Vi kommer särskilt att leta efter bevis att varje nytt förslag på ett korrekt sätt har prövats mot subsidiaritets - och proportionalitetsprinciperna , och vi kommer att leta efter sektorsspecifika debatter i Europaparlamentets egna specialiserade utskott . </s>
<s snum=175> Denna riktlinje är huvudsakligen skyddet av gemenskapens ekonomiska intressen . </s>
<s snum=176> Vi håller med er om att vi behöver ett regelbaserat handelssystem . </s>
<s snum=177> Detta är ett mycket bra exempel , men vad hände med de övriga fem ? </s>
<s snum=178> Vi krävde att kommissionen i förekommande fall lägger fram ett ändringsförslag . </s>
<s snum=179> Jag ber er därför stödja ändringsförslag 29 och 18 . </s>
<s snum=180> Det är inte heller säkert att den tredje världen sammantaget gynnas av att man förbjuder tillsatserna av andra vegetabiliska fetter . </s>
<s snum=181> Det är vad konsumenten begär . </s>
<s snum=182> Herr talman , ärade kollegor ! Jag instämmer till fullo med Luis Queirós uttalande och vilja att ytterligare tillföra debatten något . </s>
<s snum=183> Resolutionen innehåller inte mycket i den vägen , men parlamentet har redan vid minst tre tillfällen haft möjlighet att säga vad det väntade sig av en stadga om grundläggande rättigheter . </s>
<s snum=184> Vi skulle önska att den regeringskonferens som nu inleder sitt arbete hela tiden håller i minnet den viktiga regeln om respekt för de nationella demokratierna . </s>
<s snum=185> Som alla vet bör detta enligt Europaparlamentets uppfattning utgöra ett steg på vägen mot att skapa en konstitution för unionen . </s>
<s snum=186> Vi tillhör dessutom ett beprövat parti när det gäller kampen för demokrati , och vi har alltid menat att försvaret av de mänskliga rättigheterna är det absolut viktigaste . </s>
<s snum=187> Vår grupp hoppas dessutom att en nedtecknad lista över de europeiska grundläggande rättigheterna kommer att ge det europeiska integrationsvärdet ett starkare rättsligt etiskt fundament och kunna bidra till mer öppenhet och klarhet för medborgaren . </s>
<s snum=188> Det jag inte helt förstod var när han talade om andra åtgärder , då det var nödvändigt att få den gemensamma marknaden att fungera . </s>
<s snum=189> Jag vill höra er åsikt , herr kommissionär : Har ni för avsikt att vidta några åtgärder för att ekonomiskt , ekologiskt och kulturellt återställa de drabbade regionerna ? </s>
<s snum=190> Jag är övertygad om , herr kommissionär , att budgetutskottet kommer att läsa dessa uppgifter med tillfredsställelse när det får dem . </s>
<s snum=191> Eftersom ni ställer frågan kan jag säga att det land som har opponerat sig är Frankrike . </s>
<s snum=192> EU lagstiftar idag för att främja rörligheten och trafiksäkerheten . </s>
